module test #(
    
) (
    ports
);
    
endmodule